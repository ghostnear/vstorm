module vstorm

// Used to initialise the window
pub struct StormWindowConfig {
	title string
}

// Used to initialise the framework
pub struct StormConfig {
	winconfig StormWindowConfig
}
